../Simulations/Star.asc
V1 N008 0 PULSE(0 3.3 0 2e-9 1.5e-9 0.8e-8 2e-8)
R1 N004 N008 14
C1 N004 0 20e-12
R2 N005 N004 {R1}
T1 N005 0 N001 0 Td={L1} Z0={Z1}
T2 N002 0 N003 0 Td={L} Z0={Z}
T3 N006 0 N007 0 Td={L} Z0={Z}
T4 N009 0 N010 0 Td={L} Z0={Z}
R3 N002 N001 {R}
R4 N006 N001 {R}
R5 N009 N001 {R}
R6 N003 0 1e6
R7 N007 0 1e6
R8 N010 0 1e6
.tran 4e-8
.params R1 = 50.0
.params R = 50.0
.params Z1 = 50.0
.params Z = 50.0
.params L1 = 0.3537981505124526n
.params L = 0.3537981505124526n
.backanno.end