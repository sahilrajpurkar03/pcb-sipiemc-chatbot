
V1 N007 0 PULSE(0 1.5 0 2e-9 1.5e-9 0.875e-8 2e-8)
R1 N002 N007 31
C1 N002 0 20e-12
T1 N002 0 N003 0 Td={TD1} Z0={Z}
T3 N003 0 N004 0 Td={TD2} Z0={Z}
T4 N003 0 N008 0 Td={TD5} Z0={Z}
R8 N008 0 1e6
T2 N004 0 N009 0 Td={TD5} Z0={Z}
R2 N009 0 1e6
T5 N004 0 N005 0 Td={TD3} Z0={Z}
T6 N005 0 N006 0 Td={TD4} Z0={Z}
T7 N005 0 N010 0 Td={TD5} Z0={Z}
R3 N010 0 1e6
V2 N001 0 0.75
R4 N001 N006 {RT}
.tran 4e-8
.params RT = 1.0
.params L1 = 0.7075963010249052n
.params L2 = 0.7075963010249052n
.params L3 = 0.7075963010249052n
.params L4 = 0.7075963010249052n
.params L5 = 0.7075963010249052n
.params Z = 50.0
.backanno.end